------------------------------------------------------------
-- Neander - Modulo de Memoria
------------------------------------------------------------
