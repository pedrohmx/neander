------------------------------------------------------------
-- Neander - Modulo de Controle
------------------------------------------------------------
