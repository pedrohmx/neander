------------------------------------------------------------
--	Neander - Modulo de ULA
------------------------------------------------------------
--	Componentes
--		reg AC
--		reg FLAGS
--		ULA
------------------------------------------------------------
